library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use 


entity A6_PJH_KJW is
    Port ( A : in  STD_LOGIC;
           B : in  STD_LOGIC;
           Seg_3 : out  STD_LOGIC;
           Seg_2 : out  STD_LOGIC;
           Seg_1 : out  STD_LOGIC);
end A6_PJH_KJW;

architecture Behavioral of A6_PJH_KJW is

begin


end Behavioral;

