library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_bit.all;

entity BCD_Adder_6_KJW_PJH is
    Port ( X : in unsigned(7 downto 0);
           Y : in unsigned(7 downto 0);
           Z : out unsigned(11 downto 0));
end BCD_Adder_6_KJW_PJH;

architecture Behavioral of BCD_Adder_6_KJW_PJH is

begin


end Behavioral;

